module ALU_4
(   input [2:0]en,
    input [3:0]a,
    input [3:0]b,
    output [3:0]result,
    output zero,
    output carry,
    output overflow,
    output flag
);
endmodule