module ysyx_22050019_EX_MEM (

);
endmodule