module top(
    input[1:0] sw , 
    output ledr
);

    assign c = a & b;

/*
initial begin 
    $display("Hello World"); 
    //$finish; 
end
*/
endmodule
