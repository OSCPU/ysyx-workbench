module ysyx_22050019_ID_EX (

);
endmodule