module ysyx_22050019_MEM_WB (

);
endmodule