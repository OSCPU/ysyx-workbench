module example();
endmodule
