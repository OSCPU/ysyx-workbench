module top(
  input [3:0] a,
  input [1:0] s,
  output y
);
mux41 mux41_0(
  .a(a),
  .s(s),
  .y(y)
);






endmodule
