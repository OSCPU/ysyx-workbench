module ysyx_22050019_IF_ID (

);
endmodule