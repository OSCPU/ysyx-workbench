module top(
  input a,
  input b,
  output f
);
  assign f = 0;
endmodule
