module top(
  input a,
  input b,
  output f
);
  assign f = 1;
endmodule
